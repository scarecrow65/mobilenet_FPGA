module relu6 (
    input  wire signed [31:0] data_in,
    output wire signed [31:0] data_out
);

endmodule