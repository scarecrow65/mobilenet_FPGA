module fold_controller (
    input  wire clk,
    input  wire rst_n,

    input  wire start,
    output wire fold_done,
    output wire [7:0] fold_index
);

endmodule