module tile_controller (
    input  wire clk,
    input  wire rst_n,
    input  wire start,

    output wire load_tile,
    output wire compute_tile,
    output wire store_tile,

    output wire done
);

endmodule